`timescale 1ns/1ps

module cpu #(
  parameter integer XLEN      = 32,
  parameter integer REG_NUM   = 32,
  parameter integer ADDR_SIZE = 5,
  parameter integer PC_BITS   = 12,
  parameter [PC_BITS-1:0] RESET_PC = {PC_BITS{1'b0}}
)(
  input  wire clk,
  input  wire rst
);

  // ===== Program Counter wires =====
  wire [PC_BITS-1:0] F_pc;            // current PC (Fetch stage)
  wire [PC_BITS-1:0] pc_plus_1 = F_pc + {{(PC_BITS-1){1'b0}}, 1'b1};
<<<<<<< HEAD
=======
    // NEW: Extend PC+1 to XLEN for writing to the Register File
  wire [XLEN-1:0] pc_plus_1_ext = {{ (XLEN-PC_BITS){1'b0} }, pc_plus_1};
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)

  // ===== Instruction fetch output =====
  wire [XLEN-1:0] F_inst;             // fetched instruction

  // Hazard_unit
  wire        stall_D;

  // Branch Predictor
  wire       F_BP_taken;        
  wire [PC_BITS-1:0] F_BP_target_pc; 





  // ===== ALU output wires =====
  wire [XLEN-1:0]  EX_alu_out;
  wire             EX_taken;

  // ===== PC Register =====
  pc #(
    .PCLEN(PC_BITS),
    .RESET_PC(RESET_PC)
  ) u_pc (
    .clk       (clk),
    .rst       (rst),
    .EX_taken  (EX_taken),
    .EX_alt_pc (EX_alu_out[PC_BITS-1:0]),
    .F_BP_target_pc(F_BP_target_pc),
    .stall_D   (stall_D),
    .F_pc      (F_pc)
  );


  

  // ===== I-Cache <-> Instruction Memory wires =====
  wire        Ic_mem_req;
  wire [9:0]  Ic_mem_addr;
  wire [127:0] F_mem_inst;
  wire        F_mem_valid;
  wire        F_stall;      // from I-cache to your F-stage control

  // ===== I-Cache =====
  icache u_icache (
    .clk       (clk),
    .rst       (rst),

    .F_pc        (F_pc),        // PC from F stage

    .F_mem_inst  (F_mem_inst),  // data from instruction memory
    .F_mem_valid (F_mem_valid), // valid from instruction memory

    .Ic_mem_req   (Ic_mem_req),   // request to instruction memory
    .Ic_mem_addr  (Ic_mem_addr),  // address to instruction memory

    .F_inst      (F_inst),      // instruction to F stage
    .F_stall     (F_stall)      // stall signal to F-stage/pipeline
  );

 




 
  wire [XLEN-1:0]    D_inst;
  wire [PC_BITS-1:0] D_pc;
  wire               D_BP_taken;
  wire [PC_BITS-1:0] D_BP_target_pc;
<<<<<<< HEAD
=======
  wire [XLEN-1:0]    D_link_addr; // PC+1 (extended)

>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)

  f_to_d_reg #(
    .XLEN(XLEN),
    .PC_BITS(PC_BITS)
  ) u_f2d (
    .clk      (clk),
    .rst      (rst),
    .F_pc     (F_pc),
    .F_inst   (F_inst),
    .F_BP_taken(F_BP_taken),
    .F_BP_target_pc(F_BP_target_pc),
<<<<<<< HEAD
=======
    .F_link_addr (pc_plus_1_ext), // Input

>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)
    .stall_D  (stall_D),
    .MEM_stall (MEM_stall),
    .EX_taken (EX_taken),
    .D_pc     (D_pc),
    .D_inst   (D_inst),
    .D_BP_taken(D_BP_taken),
<<<<<<< HEAD
    .D_BP_target_pc(D_BP_target_pc)
=======
    .D_BP_target_pc(D_BP_target_pc),
    .D_link_addr (D_link_addr) // Output

>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)
   
  );


  //Decoder 

  wire [5:0]        D_opc;
  wire [4:0]        D_ra;
  wire [4:0]        D_rb;
  wire [4:0]        D_rd;
  wire [10:0]       D_imd;
  wire              D_we;
  wire [3:0]        D_alu_op;       // 4-bit ALU op
  wire              D_ld;
  wire              D_str;
  wire              D_brn;
  wire              D_addi;
  wire              D_mul;
  wire              D_byt;
<<<<<<< HEAD
=======
  wire              D_jmp;
  wire              D_link_we;
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)

  decode #(
        .XLEN(XLEN)
  ) u_decode (
    .clk      (clk),
    .D_inst   (D_inst),
    .D_opc    (D_opc),
    .D_ra     (D_ra),
    .D_rb     (D_rb),
    .D_rd     (D_rd),
    .D_imd    (D_imd),
    .D_we     (D_we),
    .D_alu_op (D_alu_op),
    .D_ld     (D_ld),
    .D_str    (D_str),
    .D_byt    (D_byt),
    .D_brn    (D_brn),
    .D_addi   (D_addi),
    .D_mul    (D_mul),
<<<<<<< HEAD
    .D_jmp    (D_jmp)
=======
    .D_jmp    (D_jmp),
    .D_link_we(D_link_we)
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)
  );

  // ----- Hazard unit wires -----
  wire [1:0]  EX_D_bp;
  wire [1:0]  MEM_D_bp;
  wire [1:0]  WB_D_bp;

  // ----- Hazard unit instance -----
  Hazard_unit #(
    .XLEN(XLEN),
    .ADDR_SIZE(ADDR_SIZE)   // use reg address size, not PC bits
  ) u_Hazard_unit (
    .clk      (clk),
    .rst      (rst),
    // Decode stage
   

    .D_ra      (D_ra),
    .D_rb      (D_rb),
    .D_rd      (D_rd),
    
    

    // EX stage
    .EX_alu_out(EX_alu_out),  // (not used for detection but fine to pass)
    .EX_rd     (EX_rd),
    .EX_we     (EX_we),
    .EX_ld     (EX_ld),
    .EX_mul     (EX_mul),

    // MEM stage
    .MEM_rd    (MEM_rd),
    .MEM_we    (MEM_we),

    // WB stage
    .WB_rd     (WB_rd),
    .WB_we     (WB_we),

    // Outputs
    .stall_D   (stall_D),
    .EX_D_bp   (EX_D_bp),     // {ra, rb}
    .MEM_D_bp  (MEM_D_bp),    // {ra, rb}
    .WB_D_bp   (WB_D_bp)      // {ra, rb}
  );

  //Regfile 
  
                                    
  wire [XLEN-1:0]      D_a;      // value of raddr1
  wire [XLEN-1:0]      D_b;       // value of raddr2
  wire [XLEN-1:0]      D_a2;       // value of raddr2
  wire [XLEN-1:0]      D_b2;       // value of raddr2


<<<<<<< HEAD
=======

>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)
  regfile #(
    .XLEN(XLEN),
    .REG_NUM(REG_NUM),
    .ADDR_SIZE(ADDR_SIZE)
  ) u_regfile (
    // From Decode
    .clk        (clk),
    .D_ra       (D_ra),      // first register to read
    .D_rb       (D_rb),      // second register to read
    .D_imd      (D_imd),
    .D_pc       (D_pc),
    .D_ld       (D_ld),
    .D_str      (D_str),
    .D_brn      (D_brn),
    .D_addi     (D_addi),
    .D_jmp      (D_jmp),
    .D_mul      (D_mul),
<<<<<<< HEAD

=======
    .D_link_we  (D_link_we),      // JALX Instruction Flag
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)
    //From Hazard_unit
    .EX_D_bp    (EX_D_bp),
    .MEM_D_bp   (MEM_D_bp),
    .WB_D_bp    (WB_D_bp),

    .EX_alu_out    (EX_alu_out),   // EX result (valid when EX_D_bp used and not a load-use)
    .MEM_data_mem  (MEM_data_mem), // data a


    // From Writeback stage
    .WB_we      (WB_we),
    .WB_rd      (WB_rd),
    .WB_data_mem(WB_data_mem),
<<<<<<< HEAD
=======
    .WB_link_we (WB_link_we),   // JALX Write Enable
    .WB_link_addr(WB_link_addr), // JALX Data (PC + 1)
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)


    // Outputs to Execute
    .D_a        (D_a),
    .D_b        (D_b),
    .D_a2       (D_a2),
    .D_b2       (D_b2)
  );



  // ===== D → EX pipeline register =====


  wire [XLEN-1:0]       EX_a;
  wire [XLEN-1:0]       EX_a2;
  wire [XLEN-1:0]       EX_b;
  wire [XLEN-1:0]       EX_b2;
  wire [3:0]            EX_alu_op;
  wire [4:0]            EX_rd;
  wire                  EX_ld;
  wire                  EX_str;
  wire                  EX_byt;
  wire                  EX_we;
  wire                  EX_brn;
  wire                  EX_mul;
  wire                  EX_BP_taken;
  wire [PC_BITS-1:0]    EX_BP_target_pc;
<<<<<<< HEAD
=======
  wire [XLEN-1:0]       EX_link_addr; // JALX Link Address
  wire                  EX_link_we;   // JALX Link Write Enable
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)


  d_to_ex_reg #(
    .XLEN(XLEN)
  ) u_d_to_ex_reg (
    .clk      (clk),
    .rst      (rst),

    // From Decode/Regfile (D stage)
    .D_a      (D_a),
    .D_a2     (D_a2),
    .D_b      (D_b),
    .D_b2     (D_b2),
    .D_alu_op (D_alu_op),
    .D_brn    (D_brn),
    .D_rd     (D_rd),
    .D_ld     (D_ld),
    .D_str    (D_str),
    .D_byt    (D_byt),
    .D_jmp    (D_jmp),  
    .D_we     (D_we),
    .D_mul    (D_mul),
    .D_BP_taken(D_BP_taken),
    .D_BP_target_pc(D_BP_target_pc),
<<<<<<< HEAD
=======
    .D_link_addr (D_link_addr), // Input
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)


    .stall_D  (stall_D),
    .MEM_stall (MEM_stall),
    .EX_taken (EX_taken),


    // To Execute stage (EX)
    .EX_a     (EX_a),
    .EX_a2    (EX_a2),
    .EX_b     (EX_b),
    .EX_b2    (EX_b2),
    .EX_alu_op(EX_alu_op),
    .EX_rd    (EX_rd),
    .EX_ld    (EX_ld),
    .EX_str   (EX_str),
    .EX_byt   (EX_byt),
    .EX_we    (EX_we),
    .EX_brn   (EX_brn),
    .EX_mul   (EX_mul),
    .EX_BP_taken(EX_BP_taken),
<<<<<<< HEAD
    .EX_BP_target_pc(EX_BP_target_pc)
=======
    .EX_BP_target_pc(EX_BP_target_pc),
    .EX_link_addr (EX_link_addr), // Output
    .EX_link_we   (EX_link_we)    // Output
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)
  );


 


  // ===== ALU stage =====

  wire       EX_true_taken;       // resolved direction

  alu #(
    .XLEN(XLEN)
  ) u_alu (
    .EX_a           (EX_a),
    .EX_a2          (EX_a2),
    .EX_b           (EX_b),
    .EX_b2          (EX_b2),
    .EX_alu_op      (EX_alu_op),
    .EX_brn         (EX_brn),
<<<<<<< HEAD
    .EX_jmp         (EX_jmp),
=======
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)
    .EX_BP_taken    (EX_BP_taken),
    .EX_BP_target_pc(EX_BP_target_pc),
    .EX_alu_out     (EX_alu_out),
    .EX_taken       (EX_taken),
    .EX_true_taken  (EX_true_taken)
  );



  branch_buffer #(
  ) u_branch_buffer (
    .clk             (clk),
    .rst             (rst),
    .F_pc            (F_pc),
    .EX_brn          (EX_brn),
    .F_stall         (F_stall),
    .MEM_stall       (MEM_stall),
    .EX_pc           (EX_a[PC_BITS-1:0]),
    .EX_alu_out      (EX_alu_out[PC_BITS-1:0]),
    .EX_true_taken   (EX_true_taken),
    .F_BP_target_pc  (F_BP_target_pc),
    .F_BP_taken      (F_BP_taken)
  );



  // ===== EX → MEM pipeline register wires =====
<<<<<<< HEAD
  wire [XLEN-1:0] MEM_alu_out;
  wire             MEM_taken;
  wire [XLEN-1:0] MEM_b2;
  wire [XLEN-1:0] MEM_a2;
  wire [4:0]       MEM_rd;
  wire             MEM_we;
  wire             MEM_ld;
  wire             MEM_str;
  wire             MEM_byt;
=======
  wire [XLEN-1:0]   MEM_alu_out;
  wire              MEM_taken;
  wire [XLEN-1:0]   MEM_b2;
  wire [XLEN-1:0]   MEM_a2;
  wire [4:0]        MEM_rd;
  wire              MEM_we;
  wire              MEM_ld;
  wire              MEM_str;
  wire              MEM_byt;
  wire  [XLEN-1:0]  MEM_link_addr;
  wire              MEM_link_we;
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)


  // ===== EX → MEM pipeline register =====
  ex_to_mem_reg #(
    .XLEN(XLEN)
  ) u_ex_to_mem_reg (
    .clk        (clk),
    .rst        (rst),

    // From Execute stage (EX)
    .EX_alu_out (EX_alu_out),
    .EX_taken   (EX_taken),
    .EX_b2      (EX_b2),
    .EX_a2      (EX_a2),
    .EX_rd      (EX_rd),
    .EX_we      (EX_we),
    .EX_ld      (EX_ld),
    .EX_str     (EX_str),
    .EX_byt     (EX_byt),
    .MEM_stall (MEM_stall),
<<<<<<< HEAD
=======
    .EX_link_addr (EX_link_addr), // Input
    .EX_link_we   (EX_link_we),   // Input
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)

    // To Memory stage (MEM)
    .MEM_alu_out(MEM_alu_out),
    .MEM_taken  (MEM_taken),
    .MEM_b2     (MEM_b2),
    .MEM_a2     (MEM_a2),
    .MEM_rd     (MEM_rd),
    .MEM_we     (MEM_we),
    .MEM_ld     (MEM_ld),
    .MEM_str    (MEM_str),
<<<<<<< HEAD
    .MEM_byt    (MEM_byt)
=======
    .MEM_byt    (MEM_byt),
    .MEM_link_addr (MEM_link_addr), // Input
    .MEM_link_we   (MEM_link_we)      // Input
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)
  );






  // ============ D-cache <-> backing data memory ===============
  wire             Dc_mem_req;
  wire [9:0]       Dc_mem_addr;     // 16 lines in backing memory
  wire [127:0]     MEM_data_line;
  wire             MEM_mem_valid;

  wire             Dc_wb_we;
  wire [9:0]       Dc_wb_addr;
  wire [127:0]     Dc_wb_wline;
  wire [XLEN-1:0]  MEM_data_mem;



  dcache #(
    .XLEN(XLEN)
  ) u_dcache (
    .clk         (clk),
    .rst         (rst),
    .MEM_ld      (MEM_ld),
    .MEM_str     (MEM_str),
    .MEM_byt     (MEM_byt),
    .MEM_alu_out (MEM_alu_out),
    .MEM_b2      (MEM_b2),

    // To MEM stage
    .MEM_data_mem(MEM_data_mem),
    .MEM_stall   (MEM_stall),

    // Backing memory: line read
    .Dc_mem_req   (Dc_mem_req),
    .Dc_mem_addr  (Dc_mem_addr),
    .MEM_data_line    (MEM_data_line),
    .MEM_mem_valid (MEM_mem_valid),

    // Backing memory: line write-back
    .Dc_wb_we    (Dc_wb_we),
    .Dc_wb_addr  (Dc_wb_addr),
    .Dc_wb_wline (Dc_wb_wline)

  );

    // Unified instruction + data memory
unified_mem #(
    .XLEN    (XLEN),
    .LATENCY (3)       // same latency you used before
) u_unified_mem (
    .clk  (clk),
    .rst  (rst),

    // ================== Instruction side ==================
    .Ic_mem_req  (Ic_mem_req),   // from your fetch/I-cache
    .Ic_mem_addr (Ic_mem_addr),  // line index
    .F_mem_inst  (F_mem_inst),   // 128-bit instruction line
    .F_mem_valid (F_mem_valid),

    // ====================== Data side ======================
    // Line read
    .Dc_mem_req    (Dc_mem_req),
    .Dc_mem_addr   (Dc_mem_addr),
    .MEM_data_line (MEM_data_line),
    .MEM_mem_valid (MEM_mem_valid),

    // Line write-back
    .Dc_wb_we    (Dc_wb_we),
    .Dc_wb_addr  (Dc_wb_addr),
    .Dc_wb_wline (Dc_wb_wline)
);


  
  



  // ===== MEM → WB pipeline register wires =====
  wire [XLEN-1:0]  WB_data_mem;
  wire [4:0]       WB_rd;
  wire             WB_we;
<<<<<<< HEAD

=======
  wire  [XLEN-1:0]  WB_link_addr;
  wire              WB_link_we;
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)
  // ===== MEM → WB pipeline register =====
  mem_to_wb_reg #(
    .XLEN(XLEN)
  ) u_mem_to_wb_reg (
    .clk         (clk),
    .rst         (rst),

    // From Memory stage (MEM)
    .MEM_data_mem(MEM_data_mem),
    .MEM_rd      (MEM_rd),
    .MEM_we      (MEM_we),
<<<<<<< HEAD

    // To Writeback stage (WB)
    .WB_data_mem (WB_data_mem),
    .WB_rd       (WB_rd),
    .WB_we       (WB_we)
=======
    .MEM_link_addr (D_link_addr), // Input
    .MEM_link_we   (D_link_we),      // Input
    // To Writeback stage (WB)
    .WB_data_mem (WB_data_mem),
    .WB_rd       (WB_rd),
    .WB_we       (WB_we),
    .WB_link_addr (WB_link_addr), // Output
    .WB_link_we   (WB_link_we)    // Output
>>>>>>> 0a5a1c4 (JALX with wrong Opcode instruction)
  );
  





 

endmodule
